/*
    
    Yves Acremann, 22.2.2021
*/

// verilator lint_off IMPLICITSTATIC
// The internally used types for the calculations:
// We use two additional bits internally in order to avoid overflows
// and for more precision.
typedef logic signed [17:0] signal_t;

// Caution: angles have two additional bits internally as we need a sign
// and a bit more precision!
// Scaling of the angle: Q2.(numOfBitsAngle-1) with 1.0 corresponding to pi.
// (for example: format: Q2.16; pi corresponds to "010000000000000000")
typedef logic signed [17:0] angle_t;

// struct containing the rotation state as well as the sign
// flip of the cosinus
typedef struct packed
{
    signal_t x;
    signal_t y;
    angle_t  z;
    logic    cos_sign;
} rot_state_t;
    

// the atan lookup table (generated by tableGen.py)
parameter angle_t atan_lut[16] = '{
    18'd16384,
    18'd9672,
    18'd5110,
    18'd2594,
    18'd1302,
    18'd652,
    18'd326,
    18'd163,
    18'd81,
    18'd41,
    18'd20,
    18'd10,
    18'd5,
    18'd3,
    18'd1,
    18'd1
};
    
/**
  The Cordic algorithm implemented as a finite state machine
**/
module CORDIC(
    input logic                 clk,
    input logic                 reset,
    input logic                 tick,    // only run if 1

    input logic unsigned[15:0]  angle,   // scaled to [0..2pi[

    input logic  signed[15:0]   x_i,     // input for mixing

    output logic signed[15:0]   x_o,     // output: cos
    output logic signed[15:0]   y_o      // output: sin
    );
    
    
    
    // the states of the FSM
    typedef enum logic [1:0] {
        IDLE,
        ITERATE,
        FINISH
    } state_t;
    
    // The signals for the iterations
    rot_state_t rot_state, next_rot_state;
    
    // the state of the FSM
    state_t  state, next_state;
    logic unsigned [3:0] iteration, next_iteration;
    

    // signals needed to store the result
    logic store_result;
    //logic signed [15:0] result_x, result_y;
    rot_state_t result;
    
    
    // the Cordic state machine: transition function
    always_comb 
    begin
        // default: do nothing
        next_state = state;
        next_iteration = iteration;
        next_rot_state = rot_state;
        store_result = 0;
        
        
        case(state)
            IDLE: 
            begin
                if (tick == 1) begin
                    // prepare the rotation vector
                    next_rot_state = PrepareRotationState(angle, x_i);
                    // prepare to iterate
                    next_iteration = 4'd0;
                    next_state = ITERATE;
                end // if tick
            end // IDLE
            
            
            ITERATE: // the actual Cordic iterations:
            begin
                next_rot_state = Rotate(rot_state, iteration);
                next_iteration = iteration + 4'd1;
                if (iteration == 15) next_state = FINISH;
            end //ITERATE
            
            FINISH:
            begin
                store_result = 1;
                next_state = IDLE; 
            end // FINISH
            
            default: next_state = IDLE; 
        endcase
    end // always_comb
    
    
    // flipflops of the FSM:
    always_ff @(posedge clk)
    begin
        if (reset == 1) begin
            state <= IDLE;
            iteration <= 4'd0;
            rot_state <= 0;
				result <= 0;
        end else begin
            state <= next_state;
            iteration <= next_iteration;
            rot_state <= next_rot_state;
				// store the result when done
				if (store_result == 1)
					result <= next_rot_state;
        end // if
    end //always_ff
    
    // convert back to 16 bits and flip the sign for the cos
    assign x_o = (result.cos_sign == 1)? 16'(-result.x >>> 2) : 16'(result.x >>> 2);
    assign y_o = 16'(result.y >>> 2);
    
endmodule // CordicFSM

/**
  Perform one rotation of the Cordic algorithm and pass on the cos_sign
 **/
function rot_state_t Rotate(
    input rot_state_t to_rotate,           // the rotation state input
    input logic unsigned [3:0] iteration   // the iteration number
    );
    
    rot_state_t result;
    // pass on the cos sign:
    result.cos_sign = to_rotate.cos_sign;
    // perform the rotation and calculate the new error for the angle:
    if (to_rotate.z > 0)
        begin
            result.x = to_rotate.x - (to_rotate.y >>> iteration);
            result.y = to_rotate.y + (to_rotate.x >>> iteration);
            result.z = to_rotate.z - atan_lut[iteration];
        end else begin
            result.x = to_rotate.x + (to_rotate.y >>> iteration);
            result.y = to_rotate.y - (to_rotate.x >>> iteration);
            result.z = to_rotate.z + atan_lut[iteration];
        end //if
        
        Rotate = result;
endfunction




/**
  Preparation at the beginning:
  * Conversion to 18 bits
  * Mapping of the angle to [-pi, pi]
  * Check if the sign of the cos output needs to be flipped
**/
function rot_state_t PrepareRotationState(
        input logic unsigned [15:0] angle,         // the angle
        input logic signed   [15:0] x_i            // input for mixing
    );
    
    
    // in this unit system, pi is just the maximum integer value / 2 
    // (and we use a signed value so the first bit is the sign!).

    
    parameter PiInt = (18'sd1 <<< 16);
    parameter PiHalfInt = PiInt >> 1;
    parameter PiThreeHalfInt = PiInt+PiHalfInt;
    
    // we use one additional bit to avoid overflows
    // (and one additional bit for better precision)
    angle_t angle_signed;
    rot_state_t rot_state;
    rot_state.x = (18'(x_i)) << 1;
    rot_state.y = 0;
    
    angle_signed = (signed'(18'(angle))) << 1;
    // determine the angle mapped to [-pi/2 .. pi/2] as well as if
    // the sign of the cos needs to be flipped.
    rot_state.cos_sign = 0;
    if ((angle_signed > PiHalfInt) & (angle_signed < PiThreeHalfInt))
        rot_state.cos_sign = 1;
        
        
    // map the angle
    if (angle_signed < PiHalfInt)
        rot_state.z = angle_signed;
    else
        if (angle_signed < PiThreeHalfInt)
            rot_state.z = PiInt-angle_signed;
        else
          // caution: This is intentional in order to avoid overflows!
          // (2pi does not fit in the signal!)
          rot_state.z = (angle_signed - PiInt) - PiInt;
        
    PrepareRotationState = rot_state;
endfunction // PrepareRotationState

// verilator lint_on IMPLICITSTATIC